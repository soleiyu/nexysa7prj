//Japari 1

module japari1
(
	input	wire  [9:0]		count,  
	output wire [15:0]  	outv
);

	reg [15:0] notes [1023:0];
	assign outv = notes[count];

	initial
	begin
	//Intro
	notes[10] <= {8'd4, 8'd49};
	notes[11] <= {8'd8, 8'd45};
	notes[12] <= {8'd4, 8'd40};
	notes[13] <= {8'd8, 8'd52};
	notes[14] <= {8'd16, 8'd49};
	
	notes[15] <= {8'd2, 8'd57};
	notes[16] <= {8'd2, 8'd56};
	notes[17] <= {8'd2, 8'd57};
	notes[18] <= {8'd4, 8'd59};
	notes[19] <= {8'd2, 8'd57};
	notes[20] <= {8'd2, 8'd59};
	notes[21] <= {8'd4, 8'd61};
	notes[22] <= {8'd2, 8'd62};
	notes[23] <= {8'd2, 8'd63};
	notes[24] <= {8'd4, 8'd64};
	notes[25] <= {8'd2, 8'd61};
	notes[26] <= {8'd2, 8'd59};
	notes[27] <= {8'd2, 8'd57};
	
	notes[28] <= {8'd4, 8'd57};
	notes[29] <= {8'd4, 8'd66};
	notes[30] <= {8'd4, 8'd64};
	notes[31] <= {8'd4, 8'd57};
	notes[32] <= {8'd4, 8'd54};
	notes[33] <= {8'd4, 8'd62};
	notes[34] <= {8'd4, 8'd61};
	notes[35] <= {8'd4, 8'd59};
	notes[36] <= {8'd4, 8'd57};
	notes[37] <= {8'd12, 8'd0};
	
	notes[38] <= {8'd32, 8'd0};
	notes[39] <= {8'd8, 8'd33};
	notes[40] <= {8'd4, 8'd76};
	notes[41] <= {8'd4, 8'd0};
	
	//Amero
	notes[42] <= {8'd2, 8'd40};
	notes[43] <= {8'd2, 8'd45};
	notes[44] <= {8'd2, 8'd48};
	notes[45] <= {8'd2, 8'd45};
	notes[46] <= {8'd3, 8'd48};
	notes[47] <= {8'd1, 8'd45};
	notes[48] <= {8'd2, 8'd0};
	notes[49] <= {8'd4, 8'd48};
	notes[50] <= {8'd2, 8'd50};
	notes[51] <= {8'd2, 8'd50};
	notes[52] <= {8'd2, 8'd48};
	notes[53] <= {8'd3, 8'd50};
	notes[54] <= {8'd3, 8'd51};
	notes[55] <= {8'd2, 8'd50};
	notes[56] <= {8'd2, 8'd48};
	notes[57] <= {8'd2, 8'd45};
	notes[58] <= {8'd2, 8'd43};
	notes[59] <= {8'd6, 8'd45};
	notes[60] <= {8'd4, 8'd0};
	
	notes[61] <= {8'd2, 8'd60};
	notes[62] <= {8'd2, 8'd57};
	notes[63] <= {8'd2, 8'd55};
	notes[64] <= {8'd6, 8'd57};
	notes[65] <= {8'd4, 8'd0};
	
	notes[66] <= {8'd2, 8'd40};
	notes[67] <= {8'd2, 8'd45};
	notes[68] <= {8'd2, 8'd48};
	notes[69] <= {8'd2, 8'd45};
	notes[70] <= {8'd3, 8'd48};
	notes[71] <= {8'd1, 8'd45};
	notes[72] <= {8'd2, 8'd0};
	notes[73] <= {8'd4, 8'd48};
	notes[74] <= {8'd2, 8'd50};
	notes[75] <= {8'd2, 8'd50};
	notes[76] <= {8'd2, 8'd48};
	notes[77] <= {8'd3, 8'd50};
	notes[78] <= {8'd3, 8'd51};
	notes[79] <= {8'd2, 8'd50};
	notes[80] <= {8'd2, 8'd48};
	notes[81] <= {8'd2, 8'd45};
	notes[82] <= {8'd2, 8'd43};
	notes[83] <= {8'd6, 8'd45};
	notes[84] <= {8'd4, 8'd0};
	
	notes[85] <= {8'd4, 8'd38};
	notes[86] <= {8'd4, 8'd39};
	notes[87] <= {8'd8, 8'd40};
	
	//Bmero
	notes[88] <= {8'd2, 8'd49};
	notes[89] <= {8'd2, 8'd49};
	notes[90] <= {8'd2, 8'd49};
	notes[91] <= {8'd2, 8'd49};
	notes[92] <= {8'd2, 8'd49};
	notes[93] <= {8'd2, 8'd54};
	notes[94] <= {8'd4, 8'd49};
	
	notes[95] <= {8'd2, 8'd48};
	notes[96] <= {8'd2, 8'd48};
	notes[97] <= {8'd2, 8'd47};
	notes[98] <= {8'd2, 8'd47};
	notes[99] <= {8'd2, 8'd45};
	notes[100] <= {8'd2, 8'd45};
	notes[101] <= {8'd4, 8'd47};
	
	notes[102] <= {8'd2, 8'd47};
	notes[103] <= {8'd2, 8'd47};
	notes[104] <= {8'd2, 8'd47};
	notes[105] <= {8'd2, 8'd47};
	notes[106] <= {8'd4, 8'd52};
	notes[107] <= {8'd2, 8'd47};
	notes[108] <= {8'd2, 8'd47};
	
	notes[109] <= {8'd2, 8'd0};
	notes[110] <= {8'd2, 8'd46};
	notes[111] <= {8'd2, 8'd0};
	notes[112] <= {8'd2, 8'd47};
	notes[113] <= {8'd2, 8'd0};
	notes[114] <= {8'd2, 8'd49};
	notes[115] <= {8'd2, 8'd0};
	notes[116] <= {8'd8, 8'd50};
	notes[117] <= {8'd2, 8'd42};
	notes[118] <= {8'd4, 8'd42};
	notes[119] <= {8'd4, 8'd0};
	
	notes[120] <= {8'd6, 8'd49};
	notes[121] <= {8'd2, 8'd40};
	notes[122] <= {8'd4, 8'd40};
	notes[123] <= {8'd2, 8'd0};
	notes[124] <= {8'd2, 8'd40};
	
	notes[125] <= {8'd4, 8'd41};
	notes[126] <= {8'd2, 8'd43};
	notes[127] <= {8'd4, 8'd45};
	notes[128] <= {8'd4, 8'd52};
	notes[129] <= {8'd4, 8'd49};
	notes[130] <= {8'd2, 8'd50};
	notes[131] <= {8'd2, 8'd49};
	notes[132] <= {8'd2, 8'd49};
	notes[133] <= {8'd8, 8'd47};
	
	notes[134] <= {8'd4, 8'd0};
	notes[135] <= {8'd2, 8'd59};
	notes[136] <= {8'd2, 8'd0};
	notes[137] <= {8'd2, 8'd52};
	notes[138] <= {8'd2, 8'd0};
	notes[139] <= {8'd2, 8'd64};
	notes[140] <= {8'd2, 8'd0};
	
	//Sabi
	notes[141] <= {8'd2, 8'd57};
	notes[142] <= {8'd2, 8'd56};
	notes[143] <= {8'd2, 8'd57};
	notes[144] <= {8'd4, 8'd59};
	notes[145] <= {8'd2, 8'd57};
	notes[146] <= {8'd2, 8'd59};
	notes[147] <= {8'd4, 8'd61};
	notes[148] <= {8'd2, 8'd62};
	notes[149] <= {8'd2, 8'd63};
	notes[150] <= {8'd4, 8'd64};
	notes[151] <= {8'd2, 8'd61};
	notes[152] <= {8'd2, 8'd59};
	notes[153] <= {8'd2, 8'd57};
	
	notes[154] <= {8'd4, 8'd57};
	notes[155] <= {8'd4, 8'd66};
	notes[156] <= {8'd4, 8'd64};
	notes[157] <= {8'd4, 8'd57};
	
	notes[158] <= {8'd2, 8'd62};	
	notes[159] <= {8'd2, 8'd61};
	notes[160] <= {8'd2, 8'd59};
	notes[161] <= {8'd2, 8'd57};
	notes[162] <= {8'd4, 8'd59};
	notes[163] <= {8'd4, 8'd0};
	
	notes[164] <= {8'd2, 8'd57};
	notes[165] <= {8'd2, 8'd56};
	notes[166] <= {8'd2, 8'd57};
	notes[167] <= {8'd4, 8'd59};
	notes[168] <= {8'd2, 8'd57};
	notes[169] <= {8'd2, 8'd59};
	notes[170] <= {8'd4, 8'd61};
	notes[171] <= {8'd2, 8'd62};
	notes[172] <= {8'd2, 8'd63};
	notes[173] <= {8'd4, 8'd64};
	notes[174] <= {8'd2, 8'd61};
	notes[175] <= {8'd2, 8'd59};
	notes[176] <= {8'd2, 8'd57};
	
	notes[177] <= {8'd4, 8'd57};
	notes[178] <= {8'd4, 8'd66};
	notes[179] <= {8'd4, 8'd64};
	notes[180] <= {8'd4, 8'd57};
	 
	notes[181] <= {8'd4, 8'd54};
	notes[182] <= {8'd4, 8'd62};
	notes[183] <= {8'd4, 8'd61};
	notes[184] <= {8'd4, 8'd59};
	
	notes[185] <= {8'd8, 8'd57};
	notes[186] <= {8'd2, 8'd0};
	notes[187] <= {8'd2, 8'd57};
	notes[188] <= {8'd2, 8'd57};
	notes[189] <= {8'd2, 8'd59};
 
	notes[190] <= {8'd4, 8'd60};
	notes[191] <= {8'd4, 8'd59};
	notes[192] <= {8'd4, 8'd57};
	notes[193] <= {8'd4, 8'd54};
	
	notes[194] <= {8'd3, 8'd52};
	notes[195] <= {8'd3, 8'd61};
	notes[196] <= {8'd2, 8'd61};
	notes[197] <= {8'd3, 8'd61};
	notes[198] <= {8'd3, 8'd60};
	notes[199] <= {8'd2, 8'd61};
	
	notes[200] <= {8'd6, 8'd62};
	notes[201] <= {8'd1, 8'd64};
	notes[202] <= {8'd1, 8'd62};
	notes[203] <= {8'd4, 8'd61};
	notes[204] <= {8'd2, 8'd0};
	notes[205] <= {8'd2, 8'd61};
	
	notes[206] <= {8'd4, 8'd62};
	notes[207] <= {8'd2, 8'd61};
	notes[208] <= {8'd4, 8'd57};
	notes[209] <= {8'd4, 8'd54};
	notes[210] <= {8'd14, 8'd57};
	notes[211] <= {8'd2, 8'd1};
	notes[212] <= {8'd2, 8'd61};
	
	notes[213] <= {8'd4, 8'd62};
	notes[214] <= {8'd2, 8'd61};
	notes[215] <= {8'd4, 8'd57};
	notes[216] <= {8'd4, 8'd54};
	notes[217] <= {8'd2, 8'd54};
	
	notes[218] <= {8'd4, 8'd52};
	notes[219] <= {8'd4, 8'd0};
	notes[220] <= {8'd8, 8'd59};
	
	notes[221] <= {8'd4, 8'd57};
	notes[222] <= {8'd12, 8'd0};
 
	notes[223] <= {8'd8, 8'd33};
	notes[224] <= {8'd4, 8'd76};
	notes[225] <= {8'd4, 8'd0};
	
	//Outro
	notes[226] <= {8'd2, 8'd61};
	notes[227] <= {8'd2, 8'd57};
	notes[228] <= {8'd2, 8'd54};
	notes[229] <= {8'd6, 8'd59};
	notes[230] <= {8'd4, 8'd0};
	
	notes[231] <= {8'd2, 8'd59};
	notes[232] <= {8'd2, 8'd56};
	notes[233] <= {8'd2, 8'd52};
	notes[234] <= {8'd6, 8'd57};
	notes[235] <= {8'd4, 8'd49};
	
	notes[236] <= {8'd4, 8'd50};
	notes[237] <= {8'd4, 8'd57};
	notes[238] <= {8'd2, 8'd56};
	notes[239] <= {8'd2, 8'd57};
	notes[240] <= {8'd4, 8'd56};
	
	notes[241] <= {8'd2, 8'd54};
	notes[242] <= {8'd2, 8'd52};
	notes[243] <= {8'd2, 8'd49};
	notes[244] <= {8'd6, 8'd54};
	notes[245] <= {8'd4, 8'd0};
	
	notes[246] <= {8'd2, 8'd61};
	notes[247] <= {8'd2, 8'd57};
	notes[248] <= {8'd2, 8'd54};
	notes[249] <= {8'd6, 8'd59};
	notes[250] <= {8'd4, 8'd0};
	
	notes[251] <= {8'd2, 8'd59};
	notes[252] <= {8'd2, 8'd61};
	notes[253] <= {8'd2, 8'd62};
	notes[254] <= {8'd4, 8'd61};
	notes[255] <= {8'd2, 8'd59};
	notes[256] <= {8'd4, 8'd57};
	
	notes[257] <= {8'd4, 8'd50};
	notes[258] <= {8'd4, 8'd57};
	notes[259] <= {8'd4, 8'd56};
	notes[260] <= {8'd2, 8'd57};
	notes[261] <= {8'd2, 8'd59};
	
	notes[262] <= {8'd6, 8'd59};
	notes[263] <= {8'd2, 8'd57};
	notes[264] <= {8'd4, 8'd57};
	notes[265] <= {8'd4, 8'd0};
	//
	notes[266] <= {8'd2, 8'd61};
	notes[267] <= {8'd2, 8'd57};
	notes[268] <= {8'd2, 8'd54};
	notes[269] <= {8'd6, 8'd59};
	notes[270] <= {8'd4, 8'd0};
	
	notes[271] <= {8'd2, 8'd59};
	notes[272] <= {8'd2, 8'd56};
	notes[273] <= {8'd2, 8'd52};
	notes[274] <= {8'd6, 8'd57};
	notes[275] <= {8'd4, 8'd49};
	
	notes[276] <= {8'd4, 8'd50};
	notes[277] <= {8'd4, 8'd57};
	notes[278] <= {8'd2, 8'd56};
	notes[279] <= {8'd2, 8'd57};
	notes[280] <= {8'd4, 8'd56};
	
	notes[281] <= {8'd2, 8'd54};
	notes[282] <= {8'd2, 8'd52};
	notes[283] <= {8'd2, 8'd49};
	notes[284] <= {8'd6, 8'd54};
	notes[285] <= {8'd4, 8'd0};
	
	notes[286] <= {8'd2, 8'd61};
	notes[287] <= {8'd2, 8'd57};
	notes[288] <= {8'd2, 8'd54};
	notes[289] <= {8'd6, 8'd59};
	notes[290] <= {8'd4, 8'd0};
	
	notes[291] <= {8'd2, 8'd59};
	notes[292] <= {8'd2, 8'd61};
	notes[293] <= {8'd2, 8'd62};
	notes[294] <= {8'd4, 8'd61};
	notes[295] <= {8'd2, 8'd59};
	notes[296] <= {8'd4, 8'd57};
	
	notes[297] <= {8'd4, 8'd50};
	notes[298] <= {8'd4, 8'd57};
	notes[299] <= {8'd4, 8'd56};
	notes[300] <= {8'd2, 8'd57};
	notes[301] <= {8'd2, 8'd59};
	
	notes[302] <= {8'd6, 8'd59};
	notes[303] <= {8'd2, 8'd57};
	notes[304] <= {8'd4, 8'd57};
	notes[305] <= {8'd4, 8'd0};
	
	notes[306] <= {8'd2, 8'd50};
	notes[307] <= {8'd2, 8'd0};
	notes[308] <= {8'd2, 8'd57};
	notes[309] <= {8'd2, 8'd0};
	notes[310] <= {8'd2, 8'd56};
	notes[311] <= {8'd2, 8'd0};
	notes[312] <= {8'd2, 8'd57};
	notes[313] <= {8'd4, 8'd59};
	notes[314] <= {8'd2, 8'd57};
	notes[315] <= {8'd2, 8'd59};
	notes[316] <= {8'd2, 8'd0};
	notes[317] <= {8'd4, 8'd57};
	notes[318] <= {8'd4, 8'd0};
	end
	
endmodule

module japari2
(
	input	wire  [9:0]		count,  
	output wire [15:0]  	outv
);

	reg [15:0] notes [1023:0];
	assign outv = notes[count];

	initial
	begin

	notes[10] <= {8'd4, 8'd0};
	notes[11] <= {8'd8, 8'd0};
	notes[12] <= {8'd4, 8'd0};
	notes[13] <= {8'd8, 8'd0};
	notes[14] <= {8'd16, 8'd0};
	
	notes[15] <= {8'd2, 8'd52};
	notes[16] <= {8'd4, 8'd0};
	notes[17] <= {8'd4, 8'd53};
	notes[18] <= {8'd4, 8'd0};
	notes[19] <= {8'd4, 8'd57};
	notes[20] <= {8'd4, 8'd0};
	notes[21] <= {8'd4, 8'd59};
	notes[22] <= {8'd2, 8'd0};
	notes[23] <= {8'd2, 8'd52};
	notes[24] <= {8'd2, 8'd0};
	
	notes[25] <= {8'd4, 8'd54};
	notes[26] <= {8'd4, 8'd57};
	notes[27] <= {8'd4, 8'd57};
	notes[28] <= {8'd4, 8'd52};
	
	notes[29] <= {8'd4, 8'd50};
	notes[30] <= {8'd4, 8'd0};
	notes[31] <= {8'd4, 8'd56};
	notes[32] <= {8'd4, 8'd0};
	
	notes[33] <= {8'd4, 8'd52};
	notes[34] <= {8'd12, 8'd0};
	notes[35] <= {8'd48, 8'd0};
	
	//A
	notes[36] <= {8'd2, 8'd37};
	notes[37] <= {8'd6, 8'd0};
	notes[38] <= {8'd3, 8'd43};
	notes[39] <= {8'd3, 8'd0};
	notes[40] <= {8'd4, 8'd45};
	notes[41] <= {8'd6, 8'd0};
	notes[42] <= {8'd3, 8'd47};
	notes[43] <= {8'd5, 8'd0};
	
	notes[44] <= {8'd2, 8'd45};
	notes[45] <= {8'd14, 8'd0};
	
	notes[46] <= {8'd2, 8'd57};
	notes[47] <= {8'd14, 8'd0};
	
	notes[48] <= {8'd2, 8'd37};
	notes[49] <= {8'd6, 8'd0};
	notes[50] <= {8'd3, 8'd43};
	notes[51] <= {8'd3, 8'd0};
	notes[52] <= {8'd4, 8'd45};
	notes[53] <= {8'd6, 8'd0};
	notes[54] <= {8'd8, 8'd47};
	
	notes[55] <= {8'd2, 8'd45};
	notes[56] <= {8'd14, 8'd0};
	
	notes[57] <= {8'd4, 8'd33};
	notes[58] <= {8'd4, 8'd34};
	notes[59] <= {8'd8, 8'd35};
	
	//B
	notes[60] <= {8'd2, 8'd45};
	notes[61] <= {8'd6, 8'd0};
	notes[62] <= {8'd2, 8'd42};
	notes[63] <= {8'd6, 8'd0};
	
	notes[64] <= {8'd2, 8'd45};
	notes[65] <= {8'd6, 8'd0};
	notes[66] <= {8'd2, 8'd42};
	notes[67] <= {8'd6, 8'd0};
	
	notes[68] <= {8'd2, 8'd44};
	notes[69] <= {8'd6, 8'd0};
	notes[70] <= {8'd4, 8'd40};
	notes[71] <= {8'd2, 8'd0};
	notes[72] <= {8'd2, 8'd40};
	
	notes[73] <= {8'd2, 8'd0};
	notes[74] <= {8'd2, 8'd40};
	notes[75] <= {8'd2, 8'd0};
	notes[76] <= {8'd2, 8'd40};
	notes[77] <= {8'd2, 8'd0};
	notes[78] <= {8'd2, 8'd45};
	notes[79] <= {8'd2, 8'd0};
	notes[80] <= {8'd8, 8'd42};
	notes[81] <= {8'd2, 8'd0};
	notes[82] <= {8'd4, 8'd38};
	notes[83] <= {8'd4, 8'd0};
	
	notes[84] <= {8'd6, 8'd45};
	notes[85] <= {8'd2, 8'd0};
	notes[86] <= {8'd4, 8'd37};
	notes[87] <= {8'd4, 8'd0};
	
	notes[88] <= {8'd4, 8'd36};
	notes[89] <= {8'd2, 8'd0};
	notes[90] <= {8'd4, 8'd41};
	notes[91] <= {8'd4, 8'd0};
	notes[92] <= {8'd4, 8'd45};
	notes[93] <= {8'd6, 8'd0};
	notes[94] <= {8'd8, 8'd44};
	
	notes[95] <= {8'd16, 8'd0};
	
	//Sabi
	notes[96] <= {8'd2, 8'd52};
	notes[97] <= {8'd4, 8'd52};
	notes[98] <= {8'd4, 8'd53};
	notes[99] <= {8'd4, 8'd53};
	notes[100] <= {8'd4, 8'd57};
	notes[101] <= {8'd4, 8'd57};
	notes[102] <= {8'd4, 8'd59};
	notes[103] <= {8'd2, 8'd59};
	notes[104] <= {8'd2, 8'd52};
	notes[105] <= {8'd2, 8'd52};
	
	notes[106] <= {8'd4, 8'd54};
	notes[107] <= {8'd4, 8'd57};
	notes[108] <= {8'd4, 8'd57};
	notes[109] <= {8'd4, 8'd52};
	
	notes[110] <= {8'd2, 8'd54};
	notes[111] <= {8'd6, 8'd544};
	notes[112] <= {8'd4, 8'd56};
	notes[113] <= {8'd4, 8'd0};
	
	notes[114] <= {8'd2, 8'd52};
	notes[115] <= {8'd4, 8'd52};
	notes[116] <= {8'd4, 8'd53};
	notes[117] <= {8'd4, 8'd53};
	notes[118] <= {8'd4, 8'd57};
	notes[119] <= {8'd4, 8'd57};
	notes[120] <= {8'd4, 8'd59};
	notes[121] <= {8'd2, 8'd59};
	notes[122] <= {8'd2, 8'd52};
	notes[123] <= {8'd2, 8'd52};
	
	notes[124] <= {8'd4, 8'd54};
	notes[125] <= {8'd4, 8'd57};
	notes[126] <= {8'd4, 8'd57};
	notes[127] <= {8'd4, 8'd52};
	
	notes[128] <= {8'd4, 8'd50};
	notes[129] <= {8'd4, 8'd50};
	notes[130] <= {8'd4, 8'd56};
	notes[131] <= {8'd4, 8'd56};
	
	notes[132] <= {8'd8, 8'd53};
	notes[133] <= {8'd8, 8'd0};
	
	
	notes[134] <= {8'd4, 8'd57};
	notes[135] <= {8'd4, 8'd57};
	notes[136] <= {8'd4, 8'd54};
	notes[137] <= {8'd4, 8'd54};
	
	notes[138] <= {8'd3, 8'd49};
	notes[139] <= {8'd5, 8'd0};
	notes[140] <= {8'd3, 8'd52};
	notes[141] <= {8'd5, 8'd0};
	
	notes[142] <= {8'd6, 8'd55};
	notes[143] <= {8'd2, 8'd55};
	notes[144] <= {8'd4, 8'd57};
	notes[145] <= {8'd4, 8'd57};
 
	notes[146] <= {8'd4, 8'd54};
	notes[147] <= {8'd2, 8'd54};
	notes[148] <= {8'd4, 8'd54};
	notes[149] <= {8'd4, 8'd0};
	notes[150] <= {8'd2, 8'd49};
	
	notes[151] <= {8'd4, 8'd50};
	notes[152] <= {8'd2, 8'd49};
	notes[153] <= {8'd4, 8'd45};
	notes[154] <= {8'd4, 8'd42};
	notes[155] <= {8'd2, 8'd0};
	
	notes[156] <= {8'd4, 8'd57};
	notes[157] <= {8'd2, 8'd57};
	notes[158] <= {8'd4, 8'd54};
	notes[159] <= {8'd4, 8'd54};
	notes[160] <= {8'd2, 8'd0};
	
	notes[161] <= {8'd4, 8'd47};
	notes[162] <= {8'd4, 8'd0};
	notes[163] <= {8'd8, 8'd47};
	
	notes[164] <= {8'd4, 8'd52};
	notes[165] <= {8'd12, 8'd0};
	
	notes[166] <= {8'd16, 8'd0};
	
	//outro
	notes[167] <= {8'd2, 8'd54};
	notes[168] <= {8'd2, 8'd54};
	notes[169] <= {8'd2, 8'd0};
	notes[170] <= {8'd6, 8'd56};
	notes[171] <= {8'd4, 8'd0};
	
	notes[172] <= {8'd2, 8'd56};
	notes[173] <= {8'd2, 8'd0};
	notes[174] <= {8'd2, 8'd0};
	notes[175] <= {8'd6, 8'd52};
	notes[176] <= {8'd4, 8'd45};
	
	notes[177] <= {8'd4, 8'd45};
	notes[178] <= {8'd4, 8'd45};
	notes[179] <= {8'd2, 8'd50};
	notes[180] <= {8'd2, 8'd50};
	notes[181] <= {8'd4, 8'd50};
	
	notes[182] <= {8'd2, 8'd48};
	notes[183] <= {8'd2, 8'd48};
	notes[184] <= {8'd2, 8'd0};
	notes[185] <= {8'd6, 8'd48};
	notes[186] <= {8'd4, 8'd0};
	
	notes[187] <= {8'd2, 8'd54};
	notes[188] <= {8'd2, 8'd54};
	notes[189] <= {8'd2, 8'd0};
	notes[190] <= {8'd6, 8'd56};
	notes[191] <= {8'd4, 8'd0};
	
	notes[192] <= {8'd2, 8'd56};
	notes[193] <= {8'd2, 8'd56};
	notes[194] <= {8'd2, 8'd56};
	notes[195] <= {8'd4, 8'd57};
	notes[196] <= {8'd2, 8'd0};
	notes[197] <= {8'd4, 8'd52};
	
	notes[198] <= {8'd4, 8'd47};
	notes[199] <= {8'd4, 8'd47};
	notes[200] <= {8'd4, 8'd50};
	notes[201] <= {8'd4, 8'd50};
		
	notes[202] <= {8'd6, 8'd52};
	notes[203] <= {8'd2, 8'd52};
	notes[204] <= {8'd4, 8'd52};
	notes[205] <= {8'd4, 8'd0};
	
	notes[206] <= {8'd2, 8'd54};
	notes[207] <= {8'd2, 8'd54};
	notes[208] <= {8'd2, 8'd0};
	notes[209] <= {8'd6, 8'd56};
	notes[210] <= {8'd4, 8'd0};
	
	notes[211] <= {8'd2, 8'd56};
	notes[212] <= {8'd2, 8'd0};
	notes[213] <= {8'd2, 8'd0};
	notes[214] <= {8'd6, 8'd52};
	notes[215] <= {8'd4, 8'd45};
	
	notes[216] <= {8'd4, 8'd45};
	notes[217] <= {8'd4, 8'd45};
	notes[218] <= {8'd2, 8'd50};
	notes[219] <= {8'd2, 8'd50};
	notes[220] <= {8'd4, 8'd50};
	
	notes[221] <= {8'd2, 8'd48};
	notes[222] <= {8'd2, 8'd48};
	notes[223] <= {8'd2, 8'd0};
	notes[224] <= {8'd6, 8'd48};
	notes[225] <= {8'd4, 8'd0};
	
	notes[226] <= {8'd2, 8'd54};
	notes[227] <= {8'd2, 8'd54};
	notes[228] <= {8'd2, 8'd0};
	notes[229] <= {8'd6, 8'd56};
	notes[230] <= {8'd4, 8'd0};
	
	notes[231] <= {8'd2, 8'd56};
	notes[232] <= {8'd2, 8'd56};
	notes[233] <= {8'd2, 8'd56};
	notes[234] <= {8'd4, 8'd57};
	notes[235] <= {8'd2, 8'd0};
	notes[236] <= {8'd4, 8'd52};
 
	notes[237] <= {8'd4, 8'd47};
	notes[238] <= {8'd4, 8'd47};
	notes[239] <= {8'd4, 8'd50};
	notes[240] <= {8'd4, 8'd50};
		
	notes[241] <= {8'd6, 8'd52};
	notes[242] <= {8'd2, 8'd52};
	notes[243] <= {8'd4, 8'd52};
	notes[244] <= {8'd4, 8'd0};
	
	notes[245] <= {8'd2, 8'd45};
	notes[246] <= {8'd2, 8'd0};
	notes[247] <= {8'd2, 8'd50};
	notes[248] <= {8'd2, 8'd0};
	notes[249] <= {8'd2, 8'd50};
	notes[250] <= {8'd2, 8'd0};
	notes[251] <= {8'd2, 8'd50};
	notes[252] <= {8'd4, 8'd52};
	notes[253] <= {8'd2, 8'd52};
	notes[254] <= {8'd2, 8'd52};
	notes[255] <= {8'd2, 8'd0};
	notes[256] <= {8'd4, 8'd52};
	notes[257] <= {8'd4, 8'd0};
	
	end
endmodule

module japari3
(
	input	wire  [9:0]		count,  
	output wire [15:0]  	outv
);

	reg [15:0] notes [1023:0];
	assign outv = notes[count];

	initial
	begin
	
	notes[10] <= {8'd8, 8'd0};
	notes[11] <= {8'd12, 8'd69};
	notes[12] <= {8'd12, 8'd73};
	notes[13] <= {8'd8, 8'd69};	
	
	notes[14] <= {8'd2, 8'd33};
	notes[15] <= {8'd4, 8'd0};
	notes[16] <= {8'd2, 8'd32};
	notes[17] <= {8'd6, 8'd0};
	notes[18] <= {8'd2, 8'd30};
	
	notes[19] <= {8'd2, 8'd0};
	notes[20] <= {8'd2, 8'd30};
	notes[21] <= {8'd2, 8'd29};
	notes[22] <= {8'd4, 8'd28};
	notes[23] <= {8'd2, 8'd16};
	notes[24] <= {8'd4, 8'd33};
	
	notes[25] <= {8'd2, 8'd26};
	notes[26] <= {8'd2, 8'd26};
	notes[27] <= {8'd2, 8'd38};
	notes[28] <= {8'd2, 8'd26};
	notes[29] <= {8'd2, 8'd25};
	notes[30] <= {8'd2, 8'd13};
	notes[31] <= {8'd2, 8'd25};
	notes[32] <= {8'd2, 8'd13};
	
	notes[33] <= {8'd2, 8'd23};
	notes[34] <= {8'd2, 8'd25};
	notes[35] <= {8'd2, 8'd26};
	notes[36] <= {8'd4, 8'd28};
	notes[37] <= {8'd2, 8'd30};
	notes[38] <= {8'd2, 8'd31};
	notes[39] <= {8'd2, 8'd32};
	
	//
	notes[40] <= {8'd2, 8'd21};
	notes[41] <= {8'd1, 8'd21};
	notes[42] <= {8'd1, 8'd33};
	notes[43] <= {8'd2, 8'd20};
	notes[44] <= {8'd1, 8'd20};
	notes[45] <= {8'd1, 8'd32};
	notes[46] <= {8'd2, 8'd19};
	notes[47] <= {8'd1, 8'd19};
	notes[48] <= {8'd1, 8'd31};
	notes[49] <= {8'd2, 8'd18};
	notes[50] <= {8'd1, 8'd30};
	notes[51] <= {8'd1, 8'd30};
 
	notes[52] <= {8'd2, 8'd17};
	notes[53] <= {8'd1, 8'd17};
	notes[54] <= {8'd1, 8'd29};
	notes[55] <= {8'd2, 8'd16};
	notes[56] <= {8'd1, 8'd16};
	notes[57] <= {8'd1, 8'd28};
	notes[58] <= {8'd2, 8'd15};
	notes[59] <= {8'd1, 8'd15};
	notes[60] <= {8'd1, 8'd17};
	notes[61] <= {8'd2, 8'd16};
	notes[62] <= {8'd1, 8'd16};
	notes[63] <= {8'd1, 8'd28};
	
	notes[64] <= {8'd2, 8'd21};
	notes[65] <= {8'd1, 8'd21};
	notes[66] <= {8'd1, 8'd33};
	notes[67] <= {8'd2, 8'd20};
	notes[68] <= {8'd1, 8'd20};
	notes[69] <= {8'd1, 8'd32};
	notes[70] <= {8'd2, 8'd19};
	notes[71] <= {8'd1, 8'd19};
	notes[72] <= {8'd1, 8'd31};
	notes[73] <= {8'd2, 8'd18};
	notes[74] <= {8'd1, 8'd30};
	notes[75] <= {8'd1, 8'd30};
	
	notes[76] <= {8'd2, 8'd17};
	notes[77] <= {8'd1, 8'd17};
	notes[78] <= {8'd1, 8'd29};
	notes[79] <= {8'd2, 8'd16};
	notes[80] <= {8'd1, 8'd16};
	notes[81] <= {8'd1, 8'd28};
	notes[82] <= {8'd2, 8'd15};
	notes[83] <= {8'd1, 8'd15};
	notes[84] <= {8'd1, 8'd17};
	notes[85] <= {8'd2, 8'd16};
	notes[86] <= {8'd1, 8'd16};
	notes[87] <= {8'd1, 8'd28};
	
	//A
	notes[88] <= {8'd8, 8'd33};
	//notes[88] <= {8'd6, 8'd0};
	notes[89] <= {8'd2, 8'd31};
	notes[90] <= {8'd4, 8'd0};
	notes[91] <= {8'd4, 8'd29};
	notes[92] <= {8'd6, 8'd0};
	notes[93] <= {8'd8, 8'd28};
	
	notes[94] <= {8'd2, 8'd21};
	notes[95] <= {8'd1, 8'd21};
	notes[96] <= {8'd1, 8'd33};
	notes[97] <= {8'd2, 8'd20};
	notes[98] <= {8'd1, 8'd20};
	notes[99] <= {8'd1, 8'd32};
	notes[100] <= {8'd2, 8'd19};
	notes[101] <= {8'd1, 8'd19};
	notes[102] <= {8'd1, 8'd31};
	notes[103] <= {8'd2, 8'd18};
	notes[104] <= {8'd1, 8'd30};
	notes[105] <= {8'd1, 8'd30};
	
	notes[106] <= {8'd2, 8'd17};
	notes[107] <= {8'd1, 8'd17};
	notes[108] <= {8'd1, 8'd29};
	notes[109] <= {8'd2, 8'd16};
	notes[110] <= {8'd1, 8'd16};
	notes[111] <= {8'd1, 8'd28};
	notes[112] <= {8'd2, 8'd15};
	notes[113] <= {8'd1, 8'd15};
	notes[114] <= {8'd1, 8'd17};
	notes[115] <= {8'd2, 8'd16};
	notes[116] <= {8'd1, 8'd16};
	notes[117] <= {8'd1, 8'd28};
	
	notes[118] <= {8'd6, 8'd33};
	notes[119] <= {8'd2, 8'd21};
	notes[120] <= {8'd2, 8'd31};
	notes[121] <= {8'd2, 8'd19};
	notes[122] <= {8'd2, 8'd31};
	notes[123] <= {8'd4, 8'd29};
	notes[124] <= {8'd2, 8'd17};
	notes[125] <= {8'd2, 8'd29};
	notes[126] <= {8'd2, 8'd17};
	notes[127] <= {8'd8, 8'd28};
	
	notes[128] <= {8'd2, 8'd21};
	notes[129] <= {8'd1, 8'd21};
	notes[130] <= {8'd1, 8'd33};
	notes[131] <= {8'd2, 8'd20};
	notes[132] <= {8'd1, 8'd20};
	notes[133] <= {8'd1, 8'd32};
	notes[134] <= {8'd2, 8'd19};
	notes[135] <= {8'd1, 8'd19};
	notes[136] <= {8'd1, 8'd31};
	notes[137] <= {8'd2, 8'd18};
	notes[138] <= {8'd1, 8'd30};
	notes[139] <= {8'd1, 8'd30};
	
	notes[140] <= {8'd4, 8'd26};
	notes[141] <= {8'd4, 8'd27};
	notes[142] <= {8'd4, 8'd28};
	notes[143] <= {8'd4, 8'd0};
	
	//B
	notes[144] <= {8'd6, 8'd27};
	notes[145] <= {8'd2, 8'd27};
	notes[146] <= {8'd6, 8'd37};
	notes[147] <= {8'd2, 8'd15};
	
	notes[148] <= {8'd6, 8'd26};
	notes[149] <= {8'd2, 8'd26};
	notes[150] <= {8'd6, 8'd36};
	notes[151] <= {8'd2, 8'd14};
	
	notes[152] <= {8'd6, 8'd25};
	notes[153] <= {8'd2, 8'd25};
	notes[154] <= {8'd4, 8'd35};
	notes[155] <= {8'd2, 8'd25};
	notes[156] <= {8'd2, 8'd31};
	
	notes[157] <= {8'd2, 8'd0};
	notes[158] <= {8'd2, 8'd31};
	notes[159] <= {8'd2, 8'd0};
	notes[160] <= {8'd2, 8'd31};
	notes[161] <= {8'd2, 8'd0};
	notes[162] <= {8'd2, 8'd30};
	notes[163] <= {8'd2, 8'd0};
	notes[164] <= {8'd4, 8'd23};
	notes[165] <= {8'd2, 8'd23};
	notes[166] <= {8'd2, 8'd35};
	notes[167] <= {8'd4, 8'd23};
	notes[168] <= {8'd2, 8'd11};
	notes[169] <= {8'd2, 8'd23};
	notes[170] <= {8'd2, 8'd11};
	
	notes[171] <= {8'd2, 8'd25};
	notes[172] <= {8'd2, 8'd25};
	notes[173] <= {8'd2, 8'd37};
	notes[174] <= {8'd4, 8'd25};
	notes[175] <= {8'd2, 8'd13};
	notes[176] <= {8'd2, 8'd25};
	notes[177] <= {8'd2, 8'd13};
	
	notes[178] <= {8'd2, 8'd26};
	notes[179] <= {8'd2, 8'd14};
	notes[180] <= {8'd2, 8'd26};
	notes[181] <= {8'd4, 8'd26};
	notes[182] <= {8'd2, 8'd14};
	notes[183] <= {8'd2, 8'd26};
	notes[184] <= {8'd4, 8'd28};
	notes[185] <= {8'd2, 8'd28};
	notes[186] <= {8'd2, 8'd26};
	notes[187] <= {8'd2, 8'd27};
	notes[188] <= {8'd2, 8'd28};
	notes[189] <= {8'd2, 8'd25};
	notes[190] <= {8'd2, 8'd26};
	notes[191] <= {8'd2, 8'd27};
	
	notes[192] <= {8'd2, 8'd28};
	notes[193] <= {8'd14, 8'd0};
	
	//Sabi
	notes[194] <= {8'd2, 8'd33};
	notes[195] <= {8'd2, 8'd21};
	notes[196] <= {8'd2, 8'd37};
	notes[197] <= {8'd4, 8'd32};
	notes[198] <= {8'd2, 8'd25};
	notes[199] <= {8'd2, 8'd32};
	notes[200] <= {8'd4, 8'd30};
	notes[201] <= {8'd2, 8'd30};
	notes[202] <= {8'd2, 8'd29};
	notes[203] <= {8'd4, 8'd28};
	notes[204] <= {8'd2, 8'd33};
	notes[205] <= {8'd2, 8'd21};
	notes[206] <= {8'd2, 8'd33};
	
	notes[207] <= {8'd2, 8'd26};
	notes[208] <= {8'd2, 8'd26};
	notes[209] <= {8'd2, 8'd38};
	notes[210] <= {8'd2, 8'd26};
	notes[211] <= {8'd2, 8'd25};
	notes[212] <= {8'd2, 8'd13};
	notes[213] <= {8'd2, 8'd25};
	notes[214] <= {8'd2, 8'd13};
	
	notes[215] <= {8'd2, 8'd23};
	notes[216] <= {8'd2, 8'd25};
	notes[217] <= {8'd2, 8'd26};
	notes[218] <= {8'd4, 8'd28};
	notes[219] <= {8'd2, 8'd30};
	notes[220] <= {8'd2, 8'd31};
	notes[221] <= {8'd2, 8'd32};
	
	notes[222] <= {8'd2, 8'd33};
	notes[223] <= {8'd2, 8'd21};
	notes[224] <= {8'd2, 8'd37};
	notes[225] <= {8'd4, 8'd32};
	notes[226] <= {8'd2, 8'd25};
	notes[227] <= {8'd2, 8'd32};
	notes[228] <= {8'd4, 8'd30};
	notes[229] <= {8'd2, 8'd30};
	notes[230] <= {8'd2, 8'd29};
	notes[231] <= {8'd4, 8'd28};
	notes[232] <= {8'd2, 8'd33};
	notes[233] <= {8'd2, 8'd21};
	notes[234] <= {8'd2, 8'd33};
	
	notes[235] <= {8'd2, 8'd26};
	notes[236] <= {8'd2, 8'd26};
	notes[237] <= {8'd2, 8'd38};
	notes[238] <= {8'd2, 8'd26};
	notes[239] <= {8'd2, 8'd25};
	notes[240] <= {8'd2, 8'd13};
	notes[241] <= {8'd2, 8'd25};
	notes[242] <= {8'd2, 8'd13};
	
	notes[243] <= {8'd2, 8'd23};
	notes[244] <= {8'd2, 8'd25};
	notes[245] <= {8'd2, 8'd26};
	notes[246] <= {8'd4, 8'd28};
	notes[247] <= {8'd2, 8'd16};
	notes[248] <= {8'd2, 8'd28};
	notes[249] <= {8'd2, 8'd16};
	
	//
	notes[250] <= {8'd6, 8'd29};
	notes[251] <= {8'd2, 8'd29};
	notes[252] <= {8'd6, 8'd41};
	notes[253] <= {8'd1, 8'd29};
	notes[254] <= {8'd1, 8'd17};
	
	notes[255] <= {8'd6, 8'd29};
	notes[256] <= {8'd4, 8'd41};
	notes[257] <= {8'd2, 8'd17};
	notes[258] <= {8'd2, 8'd29};
	notes[259] <= {8'd2, 8'd17};
 
	notes[260] <= {8'd6, 8'd33};
	notes[261] <= {8'd2, 8'd33};
	notes[262] <= {8'd6, 8'd45};
	notes[263] <= {8'd1, 8'd33};
	notes[264] <= {8'd1, 8'd21};
	
	notes[265] <= {8'd6, 8'd33};
	notes[266] <= {8'd4, 8'd45};
	notes[267] <= {8'd2, 8'd21};
	notes[268] <= {8'd2, 8'd33};
	notes[269] <= {8'd2, 8'd21};
	
	notes[270] <= {8'd2, 8'd23};
	notes[271] <= {8'd2, 8'd23};
	notes[272] <= {8'd2, 8'd35};
	notes[273] <= {8'd4, 8'd23};
	notes[274] <= {8'd2, 8'd11};
	notes[275] <= {8'd2, 8'd23};
	notes[276] <= {8'd2, 8'd11};
	
	notes[277] <= {8'd2, 8'd23};
	notes[278] <= {8'd2, 8'd11};
	notes[279] <= {8'd2, 8'd23};
	notes[280] <= {8'd4, 8'd23};
	notes[281] <= {8'd2, 8'd11};
	notes[282] <= {8'd2, 8'd23};
	notes[283] <= {8'd2, 8'd11};
	
	notes[284] <= {8'd2, 8'd28};
	notes[285] <= {8'd2, 8'd16};
	notes[286] <= {8'd2, 8'd28};
	notes[287] <= {8'd4, 8'd28};
	notes[288] <= {8'd2, 8'd16};
	notes[289] <= {8'd2, 8'd28};
	notes[290] <= {8'd2, 8'd16};
	
	notes[291] <= {8'd4, 8'd28};
	notes[292] <= {8'd12, 8'd0};
	
	notes[293] <= {8'd2, 8'd21};
	notes[294] <= {8'd1, 8'd21};
	notes[295] <= {8'd1, 8'd33};
	notes[296] <= {8'd2, 8'd20};
	notes[297] <= {8'd1, 8'd20};
	notes[298] <= {8'd1, 8'd32};
	notes[299] <= {8'd2, 8'd19};
	notes[300] <= {8'd1, 8'd19};
	notes[301] <= {8'd1, 8'd31};
	notes[302] <= {8'd2, 8'd18};
	notes[303] <= {8'd1, 8'd18};
	notes[304] <= {8'd1, 8'd30};
	
	notes[305] <= {8'd2, 8'd17};
	notes[306] <= {8'd1, 8'd17};
	notes[307] <= {8'd1, 8'd29};
	notes[308] <= {8'd2, 8'd16};
	notes[309] <= {8'd1, 8'd16};
	notes[310] <= {8'd1, 8'd28};
	notes[311] <= {8'd2, 8'd15};
	notes[312] <= {8'd1, 8'd15};
	notes[313] <= {8'd1, 8'd27};
	notes[314] <= {8'd2, 8'd16};
	notes[315] <= {8'd1, 8'd16};
	notes[316] <= {8'd1, 8'd28};
	
	//outro
	notes[317] <= {8'd2, 8'd26};
	notes[318] <= {8'd2, 8'd26};
	notes[319] <= {8'd2, 8'd38};
	notes[320] <= {8'd2, 8'd26};
	notes[321] <= {8'd2, 8'd28};
	notes[322] <= {8'd2, 8'd16};
	notes[323] <= {8'd2, 8'd32};
	notes[324] <= {8'd2, 8'd16};
	
	notes[325] <= {8'd2, 8'd25};
	notes[326] <= {8'd2, 8'd13};
	notes[327] <= {8'd2, 8'd25};
	notes[328] <= {8'd2, 8'd13};
	notes[329] <= {8'd2, 8'd24};
	notes[330] <= {8'd2, 8'd12};
	notes[331] <= {8'd2, 8'd24};
	notes[332] <= {8'd2, 8'd12};
	
	notes[333] <= {8'd2, 8'd23};
	notes[334] <= {8'd2, 8'd11};
	notes[335] <= {8'd2, 8'd23};
	notes[336] <= {8'd2, 8'd11};
	notes[337] <= {8'd2, 8'd28};
	notes[338] <= {8'd2, 8'd16};
	notes[339] <= {8'd2, 8'd32};
	notes[340] <= {8'd2, 8'd16};
	
	notes[341] <= {8'd2, 8'd33};
	notes[342] <= {8'd2, 8'd21};
	notes[343] <= {8'd2, 8'd37};
	notes[344] <= {8'd4, 8'd33};
	notes[345] <= {8'd2, 8'd21};
	notes[346] <= {8'd2, 8'd33};
	notes[347] <= {8'd2, 8'd21};
	
	notes[348] <= {8'd2, 8'd26};
	notes[349] <= {8'd2, 8'd26};
	notes[350] <= {8'd2, 8'd38};
	notes[351] <= {8'd2, 8'd26};
	notes[352] <= {8'd2, 8'd28};
	notes[353] <= {8'd2, 8'd16};
	notes[354] <= {8'd2, 8'd32};
	notes[355] <= {8'd2, 8'd16};
 
	notes[356] <= {8'd2, 8'd25};
	notes[357] <= {8'd2, 8'd13};
	notes[358] <= {8'd2, 8'd25};
	notes[359] <= {8'd2, 8'd13};
	notes[360] <= {8'd2, 8'd30};
	notes[361] <= {8'd2, 8'd18};
	notes[362] <= {8'd2, 8'd33};
	notes[363] <= {8'd2, 8'd18};
	
	notes[364] <= {8'd2, 8'd23};
	notes[365] <= {8'd2, 8'd11};
	notes[366] <= {8'd2, 8'd23};
	notes[367] <= {8'd2, 8'd11};
	notes[368] <= {8'd2, 8'd28};
	notes[369] <= {8'd2, 8'd16};
	notes[370] <= {8'd2, 8'd28};
	notes[371] <= {8'd2, 8'd16};
	
	notes[372] <= {8'd2, 8'd33};
	notes[373] <= {8'd2, 8'd21};
	notes[374] <= {8'd2, 8'd37};
	notes[375] <= {8'd4, 8'd33};
	notes[376] <= {8'd2, 8'd21};
	notes[377] <= {8'd2, 8'd33};
	notes[378] <= {8'd2, 8'd21};
	
	//
	notes[379] <= {8'd2, 8'd26};
	notes[380] <= {8'd2, 8'd14};
	notes[381] <= {8'd2, 8'd26};
	notes[382] <= {8'd2, 8'd14};
	notes[383] <= {8'd2, 8'd28};
	notes[384] <= {8'd2, 8'd16};
	notes[385] <= {8'd2, 8'd28};
	notes[386] <= {8'd2, 8'd16};
	
	notes[387] <= {8'd2, 8'd25};
	notes[388] <= {8'd2, 8'd13};
	notes[389] <= {8'd2, 8'd25};
	notes[390] <= {8'd2, 8'd13};
	notes[391] <= {8'd2, 8'd24};
	notes[392] <= {8'd2, 8'd12};
	notes[393] <= {8'd2, 8'd24};
	notes[394] <= {8'd2, 8'd12};
	
	notes[395] <= {8'd2, 8'd23};
	notes[396] <= {8'd2, 8'd11};
	notes[397] <= {8'd2, 8'd23};
	notes[398] <= {8'd2, 8'd11};
	notes[399] <= {8'd2, 8'd28};
	notes[400] <= {8'd2, 8'd16};
	notes[401] <= {8'd2, 8'd28};
	notes[402] <= {8'd2, 8'd16};
 
	notes[403] <= {8'd2, 8'd33};
	notes[404] <= {8'd2, 8'd21};
	notes[405] <= {8'd2, 8'd33};
	notes[406] <= {8'd2, 8'd21};
	notes[407] <= {8'd2, 8'd33};
	notes[408] <= {8'd2, 8'd21};
	notes[409] <= {8'd2, 8'd33};
	notes[410] <= {8'd2, 8'd21};
	
	notes[411] <= {8'd2, 8'd26};
	notes[412] <= {8'd2, 8'd14};
	notes[413] <= {8'd2, 8'd26};
	notes[414] <= {8'd2, 8'd14};
	notes[415] <= {8'd2, 8'd28};
	notes[416] <= {8'd2, 8'd16};
	notes[417] <= {8'd2, 8'd28};
	notes[418] <= {8'd2, 8'd16};
	
	notes[419] <= {8'd2, 8'd25};
	notes[420] <= {8'd2, 8'd13};
	notes[421] <= {8'd2, 8'd25};
	notes[422] <= {8'd2, 8'd13};
	notes[423] <= {8'd2, 8'd30};
	notes[424] <= {8'd2, 8'd18};
	notes[425] <= {8'd2, 8'd30};
	notes[426] <= {8'd2, 8'd18};
	
	notes[427] <= {8'd2, 8'd23};
	notes[428] <= {8'd2, 8'd11};
	notes[429] <= {8'd2, 8'd23};
	notes[430] <= {8'd2, 8'd11};
	notes[431] <= {8'd2, 8'd28};
	notes[432] <= {8'd2, 8'd16};
	notes[433] <= {8'd2, 8'd28};
	notes[434] <= {8'd2, 8'd16};
	
	notes[435] <= {8'd2, 8'd21};
	notes[436] <= {8'd2, 8'd21};
	notes[437] <= {8'd2, 8'd33};
	notes[438] <= {8'd4, 8'd21};
	notes[439] <= {8'd2, 8'd09};
	notes[440] <= {8'd2, 8'd21};
	notes[441] <= {8'd2, 8'd09};
	
	notes[442] <= {8'd2, 8'd23};
	notes[443] <= {8'd6, 8'd0};
	notes[444] <= {8'd2, 8'd28};
	notes[445] <= {8'd4, 8'd0};
	notes[446] <= {8'd4, 8'd21};
	notes[447] <= {8'd2, 8'd21};
	notes[448] <= {8'd2, 8'd33};
	notes[449] <= {8'd2, 8'd0};
	notes[450] <= {8'd4, 8'd21};
	notes[451] <= {8'd4, 8'd0};
 	
	end
endmodule
