module top
(
	input wire clk,
	input wire  [15:0] SW,
	output wire CA, CB, CC, CD, CE, CF, CG, DP,
	output wire [7:0] AN
);

endmodule
